`timescale 1ns/10ps
`include "mux2to1.v"

module programCounter(in, out, clk, reset);
	output [63:0] out;

	input [63:0] in;
	input clk, reset;

		


endmodule