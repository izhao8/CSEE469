`timescale 1ns/10ps

module forwardUnit(forA, forB, Rn, Rm, regRd, MEMrd, WBrd);
	output [1:0] forA, forb;
	
	input [4:0] Rn, Rm, MEMrd, WBrd;
	

endmodule