`timescale 1ns/10ps

module CPU ();
	
	
endmodule